`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:21:08 11/06/2014 
// Design Name: 
// Module Name:    Accumulator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Accumulator(
    input clk,
    input rst,
    input [7:0] freqSel,
    input [23:0] phaseIn,
    output [9:0] phaseOut
    );
//phase register
always @ (clk)
	begin
		if 
	end
endmodule
